/*decodificador BCD usando case
Nomes: Arthur Bracarense e Gustavo Assis
inputs [3:0]SW3
output display de 7 segmentos
*/


module decod (SW,HEX4);
input [3:0]SW;
output reg [0:6] HEX4;

always@(SW)
	begin 
		case(SW)
		4'b0000 : HEX4[0:6]= 7'b0000001;//0
		4'b0001 : HEX4[0:6]= 7'b1001111;//1
		4'b0010 : HEX4[0:6]= 7'b0010010;//2
		4'b0011 : HEX4[0:6]= 7'b0000110;//3
		4'b0100 : HEX4[0:6]= 7'b1001100;//4
		4'b0101 : HEX4[0:6]= 7'b0100100;//5
		4'b0110 : HEX4[0:6]= 7'b0100000;//6
		4'b0111 : HEX4[0:6]= 7'b0001111;//7
		4'b1000 : HEX4[0:6]= 7'b0000000;//8
		4'b1001 : HEX4[0:6]= 7'b0000100;//9
		default : HEX4[0:6]= 7'bxxxxxxx;//default
	endcase
end
	
endmodule
	
		